/* Lab Exercise 1
	Simplify the following functions using K-map and implement the circuit using logic gates.
		a) f(A,B,C,D) = ∑m (2,3,4,5,6,7,10,11,12,15)
*/

`timescale 1ns/1ns
`include "exercise1a.v"

module exercise1a_tb();

reg a, b, c, d;
wire f;

exercise1a test(f, a, b, c, d);
initial begin
        $dumpfile("exercise1a.vcd");
        $dumpvars(0, exercise1a_tb);
        
        a = 0; b = 0; c = 0; d = 0; #10;
        a = 0; b = 0; c = 0; d = 1; #10;
        a = 0; b = 0; c = 1; d = 0; #10;
        a = 0; b = 0; c = 1; d = 1; #10;
        a = 0; b = 1; c = 0; d = 0; #10;
        a = 0; b = 1; c = 0; d = 1; #10;
        a = 0; b = 1; c = 1; d = 0; #10;
        a = 0; b = 1; c = 1; d = 1; #10;
        a = 1; b = 0; c = 0; d = 0; #10;
        a = 1; b = 0; c = 0; d = 1; #10;
        a = 1; b = 0; c = 1; d = 0; #10;
        a = 1; b = 0; c = 1; d = 1; #10;
        a = 1; b = 1; c = 0; d = 0; #10;
        a = 1; b = 1; c = 0; d = 1; #10;
        a = 1; b = 1; c = 1; d = 0; #10;
        a = 1; b = 1; c = 1; d = 1; #10;
        
        $display("Test Complete");
end
endmodule
        
