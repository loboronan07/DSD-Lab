/* Lab Exercise 1a
	Implement the following functions using the specified multiplexers and write the Verilog code for
the same.
		a. F(a,b,c,d) = a’b + ac’ + abd’ + bc’d using 8 to 1 multiplexer.
*/

`timescale 1ns/1ns
`include "exercise1a.v"

module exercise1a_tb();

reg a, b, c, d;
wire f;

exercise1a test(a, b, c, d, f);
initial begin
        $dumpfile("exercise1a.vcd");
        $dumpvars(0, exercise1a_tb);
        
        a = 0; b = 0; c = 0; d = 0; #10;
        a = 0; b = 0; c = 0; d = 1; #10;
        a = 0; b = 0; c = 1; d = 0; #10;
        a = 0; b = 0; c = 1; d = 1; #10;
        a = 0; b = 1; c = 0; d = 0; #10;
        a = 0; b = 1; c = 0; d = 1; #10;
        a = 0; b = 1; c = 1; d = 0; #10;
        a = 0; b = 1; c = 1; d = 1; #10;
        a = 1; b = 0; c = 0; d = 0; #10;
        a = 1; b = 0; c = 0; d = 1; #10;
        a = 1; b = 0; c = 1; d = 0; #10;
        a = 1; b = 0; c = 1; d = 1; #10;
        a = 1; b = 1; c = 0; d = 0; #10;
        a = 1; b = 1; c = 0; d = 1; #10;
        a = 1; b = 1; c = 1; d = 0; #10;
        a = 1; b = 1; c = 1; d = 1; #10;
        
        $display("Test Complete");
end
endmodule


