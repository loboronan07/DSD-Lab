module exercise1i(f, a);
input a;
output f;
assign f = ~(~a);
endmodule